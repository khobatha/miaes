/* Machine-generated using Migen */
module ShiftRowInv(
	input [7:0] sm0,
	input [7:0] sm1,
	input [7:0] sm2,
	input [7:0] sm3,
	input [7:0] sm4,
	input [7:0] sm5,
	input [7:0] sm6,
	input [7:0] sm7,
	input [7:0] sm8,
	input [7:0] sm9,
	input [7:0] sm10,
	input [7:0] sm11,
	input [7:0] sm12,
	input [7:0] sm13,
	input [7:0] sm14,
	input [7:0] sm15,
	output [7:0] recovered0,
	output [7:0] recovered1,
	output [7:0] recovered2,
	output [7:0] recovered3,
	output [7:0] recovered4,
	output [7:0] recovered5,
	output [7:0] recovered6,
	output [7:0] recovered7,
	output [7:0] recovered8,
	output [7:0] recovered9,
	output [7:0] recovered10,
	output [7:0] recovered11,
	output [7:0] recovered12,
	output [7:0] recovered13,
	output [7:0] recovered14,
	output [7:0] recovered15
);


// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on
assign recovered0 = sm0;
assign recovered1 = sm1;
assign recovered2 = sm2;
assign recovered3 = sm3;
assign recovered4 = sm4;
assign recovered5 = sm5;
assign recovered6 = sm6;
assign recovered7 = sm7;
assign recovered8 = sm8;
assign recovered9 = sm9;
assign recovered10 = sm10;
assign recovered11 = sm11;
assign recovered12 = sm12;
assign recovered13 = sm13;
assign recovered14 = sm14;
assign recovered15 = sm15;

endmodule
