/* Machine-generated using Migen */
module ShiftRow(
	input [7:0] sm0,
	input [7:0] sm1,
	input [7:0] sm2,
	input [7:0] sm3,
	input [7:0] sm4,
	input [7:0] sm5,
	input [7:0] sm6,
	input [7:0] sm7,
	input [7:0] sm8,
	input [7:0] sm9,
	input [7:0] sm10,
	input [7:0] sm11,
	input [7:0] sm12,
	input [7:0] sm13,
	input [7:0] sm14,
	input [7:0] sm15,
	output [7:0] ctext0,
	output [7:0] ctext1,
	output [7:0] ctext2,
	output [7:0] ctext3,
	output [7:0] ctext4,
	output [7:0] ctext5,
	output [7:0] ctext6,
	output [7:0] ctext7,
	output [7:0] ctext8,
	output [7:0] ctext9,
	output [7:0] ctext10,
	output [7:0] ctext11,
	output [7:0] ctext12,
	output [7:0] ctext13,
	output [7:0] ctext14,
	output [7:0] ctext15
);


// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on
assign ctext0 = sm0;
assign ctext1 = sm1;
assign ctext2 = sm2;
assign ctext3 = sm3;
assign ctext4 = sm4;
assign ctext5 = sm5;
assign ctext6 = sm6;
assign ctext7 = sm7;
assign ctext8 = sm8;
assign ctext9 = sm9;
assign ctext10 = sm10;
assign ctext11 = sm11;
assign ctext12 = sm12;
assign ctext13 = sm13;
assign ctext14 = sm14;
assign ctext15 = sm15;

endmodule
