/* Machine-generated using Migen */
module AES_Dec(
	input [7:0] ctext0,
	input [7:0] ctext1,
	input [7:0] ctext2,
	input [7:0] ctext3,
	input [7:0] ctext4,
	input [7:0] ctext5,
	input [7:0] ctext6,
	input [7:0] ctext7,
	input [7:0] ctext8,
	input [7:0] ctext9,
	input [7:0] ctext10,
	input [7:0] ctext11,
	input [7:0] ctext12,
	input [7:0] ctext13,
	input [7:0] ctext14,
	input [7:0] ctext15,
	input [7:0] key0,
	input [7:0] key1,
	input [7:0] key2,
	input [7:0] key3,
	input [7:0] key4,
	input [7:0] key5,
	input [7:0] key6,
	input [7:0] key7,
	input [7:0] key8,
	input [7:0] key9,
	input [7:0] key10,
	input [7:0] key11,
	input [7:0] key12,
	input [7:0] key13,
	input [7:0] key14,
	input [7:0] key15,
	input [7:0] ptext0,
	input [7:0] ptext1,
	input [7:0] ptext2,
	input [7:0] ptext3,
	input [7:0] ptext4,
	input [7:0] ptext5,
	input [7:0] ptext6,
	input [7:0] ptext7,
	input [7:0] ptext8,
	input [7:0] ptext9,
	input [7:0] ptext10,
	input [7:0] ptext11,
	input [7:0] ptext12,
	input [7:0] ptext13,
	input [7:0] ptext14,
	input [7:0] ptext15
);

wire [7:0] temp_temp0;
wire [7:0] temp_temp1;
wire [7:0] temp_temp2;
wire [7:0] temp_temp3;
wire [7:0] temp_temp4;
wire [7:0] temp_temp5;
wire [7:0] temp_temp6;
wire [7:0] temp_temp7;
wire [7:0] temp_temp8;
wire [7:0] temp_temp9;
wire [7:0] temp_temp10;
wire [7:0] temp_temp11;
wire [7:0] temp_temp12;
wire [7:0] temp_temp13;
wire [7:0] temp_temp14;
wire [7:0] temp_temp15;
wire [7:0] temp1_temp10;
wire [7:0] temp1_temp11;
wire [7:0] temp1_temp12;
wire [7:0] temp1_temp13;
wire [7:0] temp1_temp14;
wire [7:0] temp1_temp15;
wire [7:0] temp1_temp16;
wire [7:0] temp1_temp17;
wire [7:0] temp1_temp18;
wire [7:0] temp1_temp19;
wire [7:0] temp1_temp110;
wire [7:0] temp1_temp111;
wire [7:0] temp1_temp112;
wire [7:0] temp1_temp113;
wire [7:0] temp1_temp114;
wire [7:0] temp1_temp115;
reg [7:0] temp215 = 1'd0;

// synthesis translate_off
reg dummy_s;
initial dummy_s <= 1'd0;
// synthesis translate_on
assign temp_temp0 = ptext0;
assign temp_temp1 = ptext1;
assign temp_temp2 = ptext2;
assign temp_temp3 = ptext3;
assign temp_temp4 = ptext4;
assign temp_temp5 = ptext5;
assign temp_temp6 = ptext6;
assign temp_temp7 = ptext7;
assign temp_temp8 = ptext8;
assign temp_temp9 = ptext9;
assign temp_temp10 = ptext10;
assign temp_temp11 = ptext11;
assign temp_temp12 = ptext12;
assign temp_temp13 = ptext13;
assign temp_temp14 = ptext14;
assign temp_temp15 = ptext15;
assign temp1_temp10 = ptext0;
assign temp1_temp11 = ptext1;
assign temp1_temp12 = ptext2;
assign temp1_temp13 = ptext3;
assign temp1_temp14 = ptext4;
assign temp1_temp15 = ptext5;
assign temp1_temp16 = ptext6;
assign temp1_temp17 = ptext7;
assign temp1_temp18 = ptext8;
assign temp1_temp19 = ptext9;
assign temp1_temp110 = ptext10;
assign temp1_temp111 = ptext11;
assign temp1_temp112 = ptext12;
assign temp1_temp113 = ptext13;
assign temp1_temp114 = ptext14;
assign temp1_temp115 = ptext15;

// synthesis translate_off
reg dummy_d;
// synthesis translate_on
always @(*) begin
	temp215 <= 1'd0;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
	temp215 <= ptext15;
// synthesis translate_off
	dummy_d <= dummy_s;
// synthesis translate_on
end

endmodule
